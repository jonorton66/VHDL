-------------------------------------------------------------------------------
--
-- Title       : pong
-- Design      : pong
-- Author      : Jon
-- Company     : Home
--
-------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\pong\pong\src\pong.vhd
-- Generated   : Sun Aug 25 20:58:53 2013
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {pong} architecture {pong}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity pong is
	 port(
		 pong : in STD_LOGIC
	     );
end pong;

--}} End of automatically maintained section

architecture pong of pong is
begin

	 -- enter your statements here --

end pong;
